module fullAdder()
endmodule
